module lr5_Prishchepa(
    input [3:0] D,    // 4-бітний вхідний сигнал
    input A0,         // адресний вхід 0
    input A1,         // адресний вхід 1
    input A2,         // адресний вхід 2
    output [3:0] Q0,  // 4-бітний вихідний сигнал 0
    output [3:0] Q1,  // 4-бітний вихідний сигнал 1
    output [3:0] Q2,  // 4-бітний вихідний сигнал 2
    output [3:0] Q3,  // 4-бітний вихідний сигнал 3
    output [3:0] Q4   // 4-бітний вихідний сигнал 4
);

    assign Q0 = (~A2 & ~A1 & ~A0) ? D : 4'b0000;
    assign Q1 = (~A2 & ~A1 &  A0) ? D : 4'b0000;
    assign Q2 = (~A2 &  A1 & ~A0) ? D : 4'b0000;
    assign Q3 = (~A2 &  A1 &  A0) ? D : 4'b0000;
    assign Q4 = ( A2 & ~A1 & ~A0) ? D : 4'b0000;

endmodule

